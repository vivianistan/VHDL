--Lab 6.2 
--Vivian Tan
--04/18/2016
--Implementing a state machine
--6 states


library ieee;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity SM is
	Port(rst, clk, X: in std_logic; 
		Q1, Q2, Q3, Z: out std_logic); 
end SM;

architecture archsm of sm is
	signal state, nextstate: integer range 0 to 5 := 0; 
	signal state_output: std_logic_vector(2 downto 0); 

begin
	state_output <= conv_std_logic_vectOr(state, 3); 
		Q3 <= state_output(2); 
		Q2 <= state_output(1); 
		Q1 <= state_output(0); 

	process(state, X)
	begin
		case State is
			when 0 =>
				if X = '0' then Z<= '0'; nextstate <= 4; 
				else Z <= '0'; nextstate <= 1; end if;
			when 1 =>
				if X = '0' then Z<= '0'; nextstate <= 2; 
				else Z <= '0'; nextstate <= 1; end if; 
			when 2 =>
				if X = '0' then Z<= '0'; nextstate <= 5; 
				else Z <= '0'; nextstate <= 3; end if; 
			when 3 =>
				if X = '0' then Z<= '1'; nextstate <= 2; 
				else Z <= '0'; nextstate <= 1; end if; 
			when 4 =>
				if X = '0' then Z<= '0'; nextstate <= 5; 
				else Z <= '0'; nextstate <= 1; end if; 
			when 5 =>
				if X = '0' then Z<= '0'; nextstate <= 5; 
				else Z <= '0'; nextstate <= 5; end if; 
 		end case; 
	end process; 

	process(clk, rst)
	begin
		if (rst = '0') then 
			state <= 0; 
		elsif clk'event and clk = '1' then  --rising edge
			state <= nextstate; 
		end if; 
	end process; 			
 
end archsm; 